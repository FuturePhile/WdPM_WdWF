module instruction_decoder (
  input wire [5:0] DATA,
  output wire ACC_CE,
  output wire [2:0] ALU_OP,
  output wire [1:0] RF_A,
  output wire [2:0] RF_SEL
);
  
always @(DATA) begin
  
end
  
endmodule