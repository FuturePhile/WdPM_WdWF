module top (
    
);
    
endmodule